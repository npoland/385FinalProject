LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY ControlUnit IS
  PORT(
      DIN : STD_LOGIC_VECTOR(3 DOWNTO 0);
      );

END ControlUnit;